`ifndef CACHE_PKG_SV
`define CACHE_PKG_SV
package cache_pkg;
	import uvm_pkg::*;
	`include "cache_item.svh"
	`include "cache_seq.svh"
	`include "cache_driver.svh"
	`include "monitor.svh"
	`include "scoreboard.svh"
	`include "agent.svh"
	`include "env.svh"
	`include "base_test.svh"
endpackage : cache_pkg 
`endif